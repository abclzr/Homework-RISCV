`include "defines.v"
module stage_id(
    input wire                  rst,
    input wire                  rdy,

    input wire[`InstAddrBus]    pc_i,
    input wire[`InstBus]        inst_i,

    input wire[]
);
endmodule : stage_id